
`include "rtl/config.svi"

module mr_ldst(
    input clk, rst

);

endmodule